library verilog;
use verilog.vl_types.all;
entity CLKBUFX4 is
    port(
        Y               : out    vl_logic;
        A               : in     vl_logic
    );
end CLKBUFX4;
