library verilog;
use verilog.vl_types.all;
entity DFFRHQX1 is
    port(
        Q               : out    vl_logic;
        D               : in     vl_logic;
        CK              : in     vl_logic;
        RN              : in     vl_logic
    );
end DFFRHQX1;
