library verilog;
use verilog.vl_types.all;
entity TIEHI is
    port(
        Y               : out    vl_logic
    );
end TIEHI;
