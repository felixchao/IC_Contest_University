library verilog;
use verilog.vl_types.all;
entity DLY4X4 is
    port(
        Y               : out    vl_logic;
        A               : in     vl_logic
    );
end DLY4X4;
