library verilog;
use verilog.vl_types.all;
entity udp_tlat is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end udp_tlat;
