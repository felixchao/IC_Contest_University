library verilog;
use verilog.vl_types.all;
entity INVXL is
    port(
        Y               : out    vl_logic;
        A               : in     vl_logic
    );
end INVXL;
