library verilog;
use verilog.vl_types.all;
entity tb_sv_unit is
end tb_sv_unit;
