library verilog;
use verilog.vl_types.all;
entity tb_term_sv_unit is
end tb_term_sv_unit;
