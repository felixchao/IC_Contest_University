library verilog;
use verilog.vl_types.all;
entity TIELO is
    port(
        Y               : out    vl_logic
    );
end TIELO;
