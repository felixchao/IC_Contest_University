library verilog;
use verilog.vl_types.all;
entity DLY4X1 is
    port(
        Y               : out    vl_logic;
        A               : in     vl_logic
    );
end DLY4X1;
