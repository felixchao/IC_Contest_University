library verilog;
use verilog.vl_types.all;
entity DLY1X4 is
    port(
        Y               : out    vl_logic;
        A               : in     vl_logic
    );
end DLY1X4;
