library verilog;
use verilog.vl_types.all;
entity udp_outrf is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end udp_outrf;
