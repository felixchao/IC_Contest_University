library verilog;
use verilog.vl_types.all;
entity testfixture1 is
end testfixture1;
