library verilog;
use verilog.vl_types.all;
entity testfixture is
end testfixture;
