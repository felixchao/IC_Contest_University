library verilog;
use verilog.vl_types.all;
entity tb_Queue is
end tb_Queue;
