library verilog;
use verilog.vl_types.all;
entity traffic_light_tb is
end traffic_light_tb;
